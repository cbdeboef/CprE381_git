library IEEE;
use IEEE.std_logic_1164.all;

package cpre381Custom is

    type std_logic_aoa is array (natural range <>) of std_logic_vector;

end package cpre381Custom;

package body cpre381Custom is 
   
end package body cpre381Custom;